module ram_128x32(data_in, addr, en, action, clk, data_out);
  
	input [6:0] addr;
	input [31:0] data_in;
	input en, clk, action;
	output [31:0] data_out;
	reg   [31:0]data_out;
	
	reg  aes_en;
	wire  d128;
	wire [127:0] e128_out;
  reg [127:0] e128_in;
	
	//reg [DATA_WIDTH-1:0] ram[2**ADDR_WIDTH-1:0];
	reg [31:0] ram[127:0];
	
	AES aes(aes_en, e128_in, e128_out, d128);
	
	always @ (posedge clk)
	begin
	  aes_en = 0;
	  if(en)
		  begin
		    //AES start
		    if(addr%5 == 0 && addr%10 != 0)  aes_en = 1;
		    //Write
		    if(action)  ram[addr] <= data_in;
		    //Read
		    else        data_out <= ram[addr];
		  end
	end
	
	always @ (aes_en)
	begin
	  e128_in <= {ram[addr-1],ram[addr-2],ram[addr-3],ram[addr-4]};
	end
	
	always @ (posedge clk)
	begin
	  if(d128)
	    begin
	       ram[addr+1] <= e128_out[31:0];
	       ram[addr+2] <= e128_out[63:32];
	       ram[addr+3] <= e128_out[95:64];
	       ram[addr+4] <= e128_out[127:96];
	       ram[addr+5] <= 32'hffffffff;
	     end
	end
  
endmodule

//0 0000010 讀出ram[2]
//0 0000011 讀出ram[3]