library verilog;
use verilog.vl_types.all;
entity aes_data_tb is
end aes_data_tb;
