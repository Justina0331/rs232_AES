module aes_data_tb;
  
	wire TX;
	reg  RX, clk, rst;
  
	rs232 f_rs232(TX, RX, clk, rst);
	initial begin
		rst = 1; clk = 0; RX = 1; //按下reset並將clk清0
	#20 rst = 0;  		   //放開reset
	
	
	////////////
	////128/////
	////////////
	
	
	///////////////////////
	///////寫入USER_KEY////
	//////////////////////
	///////////////////////////////////////////////
	////////////WRITE RAM[24](F1DDCEDB)/////////////
	///////////////////////////////////////////////
	///////////////////1_byte//////////////////////
	#1000 RX = 0;	      //開始02
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////2_byte//////////////////////
	#1000 RX = 0;       //開始 98(寫入ram[24])
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////3_byte//////////////////////
	#1000 RX = 0;       //開始 1111_0001
	#1000 RX = 1;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////4_byte//////////////////////
	#1000 RX = 0;       //開始 1101_1101
	#1000 RX = 1;       
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////5_byte//////////////////////
	#1000 RX = 0;       //開始 1100_1110
	#1000 RX = 0;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////6_byte//////////////////////
	#1000 RX = 0;       //開始 1101_1011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////7_byte//////////////////////
	#1000 RX = 0;       //開始 1100_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////8_byte//////////////////////
	#1000 RX = 0;       //開始 0000_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	#3000 RX = 1;
	///////////////////////////////////////////////
	////////////WRITE RAM[25](E2B79CE5)/////////////
	///////////////////////////////////////////////
	///////////////////1_byte//////////////////////
	#1000 RX = 0;	      //開始02
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////2_byte//////////////////////
	#1000 RX = 0;       //開始 99(寫入ram[25])
	#1000 RX = 1;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////3_byte//////////////////////
	#1000 RX = 0;       //開始 1110_0010
	#1000 RX = 0;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////4_byte//////////////////////
	#1000 RX = 0;       //開始 1011_0111
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////5_byte//////////////////////
	#1000 RX = 0;       //開始 1001_1100
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////6_byte//////////////////////
	#1000 RX = 0;       //開始 1110_0101
	#1000 RX = 1;       
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////7_byte//////////////////////
	#1000 RX = 0;       //開始 1100_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////8_byte//////////////////////
	#1000 RX = 0;       //開始 0000_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	#3000 RX = 1;
	///////////////////////////////////////////////
	////////////WRITE RAM[26](95A0ACEF)/////////////
	///////////////////////////////////////////////
	///////////////////1_byte//////////////////////
	#1000 RX = 0;	      //開始02
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////2_byte//////////////////////
	#1000 RX = 0;       //開始 9A(寫入ram[26])
	#1000 RX = 0;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////3_byte//////////////////////
	#1000 RX = 0;       //開始 1001_0101
	#1000 RX = 1;       
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////4_byte//////////////////////
	#1000 RX = 0;       //開始 1010_0000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////5_byte//////////////////////
	#1000 RX = 0;       //開始 1010_1100
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////6_byte//////////////////////
	#1000 RX = 0;       //開始 1110_1111
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////7_byte//////////////////////
	#1000 RX = 0;       //開始 1100_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////8_byte//////////////////////
	#1000 RX = 0;       //開始 0000_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	#3000 RX = 1;
	///////////////////////////////////////////////
	////////////WRITE RAM[27](838C8080)/////////////
	///////////////////////////////////////////////
	///////////////////1_byte//////////////////////
	#1000 RX = 0;	      //開始02
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////2_byte//////////////////////
	#1000 RX = 0;       //開始 9B(寫入ram[27])
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////3_byte//////////////////////
	#1000 RX = 0;       //開始 1000_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////4_byte//////////////////////
	#1000 RX = 0;       //開始 1000_1100
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////5_byte//////////////////////
	#1000 RX = 0;       //開始 1000_0000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////6_byte//////////////////////
	#1000 RX = 0;       //開始 1000_0000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////7_byte//////////////////////
	#1000 RX = 0;       //開始 1100_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////8_byte//////////////////////
	#1000 RX = 0;       //開始 0000_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	#3000 RX = 1;
	///////////////////////////////////////////////
	////////////WRITE RAM[28](80808080)/////////////
	///////////////////////////////////////////////
	///////////////////1_byte//////////////////////
	#1000 RX = 0;	      //開始02
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////2_byte//////////////////////
	#1000 RX = 0;       //開始 9C(寫入ram[28])
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////3_byte//////////////////////
	#1000 RX = 0;       //開始 1000_0000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////4_byte//////////////////////
	#1000 RX = 0;       //開始 1000_0000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////5_byte//////////////////////
	#1000 RX = 0;       //開始 1100_0000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////6_byte//////////////////////
	#1000 RX = 0;       //開始 1111_0111
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////7_byte//////////////////////
	#1000 RX = 0;       //開始 1100_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////8_byte//////////////////////
	#1000 RX = 0;       //開始 0000_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	#3000 RX = 1;
	///////////////////
	///////寫入DATA////
	///////////////////
	///////////////////////////////////////////////
	////////////WRITE RAM[4](11223344)/////////////
	///////////////////////////////////////////////
	///////////////////1_byte//////////////////////
	#1000 RX = 0;	      //開始02
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////2_byte//////////////////////
	#1000 RX = 0;       //開始 84(寫入ram[4])
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////3_byte//////////////////////
	#1000 RX = 0;       //開始 0001_0001
	#1000 RX = 1;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////4_byte//////////////////////
	#1000 RX = 0;       //開始 0010_0010
	#1000 RX = 0;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////5_byte//////////////////////
	#1000 RX = 0;       //開始 0011_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////6_byte//////////////////////
	#1000 RX = 0;       //開始 0100_0100
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////7_byte//////////////////////
	#1000 RX = 0;       //開始 1100_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////8_byte//////////////////////
	#1000 RX = 0;       //開始 0000_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	#3000 RX = 1;
	///////////////////////////////////////////////
	////////////WRITE RAM[5](22334455)/////////////
	///////////////////////////////////////////////
	///////////////////1_byte//////////////////////
	#1000 RX = 0;	      //開始02
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////2_byte//////////////////////
	#1000 RX = 0;       //開始 85(寫入ram[5])
	#1000 RX = 1;       
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////3_byte//////////////////////
	#1000 RX = 0;       //開始 0010_0010
	#1000 RX = 0;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////4_byte//////////////////////
	#1000 RX = 0;       //開始 0011_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////5_byte//////////////////////
	#1000 RX = 0;       //開始 0100_0100
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////6_byte//////////////////////
	#1000 RX = 0;       //開始 0101_0101
	#1000 RX = 1;       
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////7_byte//////////////////////
	#1000 RX = 0;       //開始 1100_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////8_byte//////////////////////
	#1000 RX = 0;       //開始 0000_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	#3000 RX = 1;
	///////////////////////////////////////////////
	////////////WRITE RAM[6](33445566)/////////////
	///////////////////////////////////////////////
	///////////////////1_byte//////////////////////
	#1000 RX = 0;	      //開始02
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////2_byte//////////////////////
	#1000 RX = 0;       //開始 86(寫入ram[6])
	#1000 RX = 0;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////3_byte//////////////////////
	#1000 RX = 0;       //開始 0011_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////4_byte//////////////////////
	#1000 RX = 0;       //開始 0100_0100
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////5_byte//////////////////////
	#1000 RX = 0;       //開始 0101_0101
	#1000 RX = 1;       
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////6_byte//////////////////////
	#1000 RX = 0;       //開始 0110_0110
	#1000 RX = 0;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////7_byte//////////////////////
	#1000 RX = 0;       //開始 1100_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////8_byte//////////////////////
	#1000 RX = 0;       //開始 0000_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	#3000 RX = 1;
	///////////////////////////////////////////////
	////////////WRITE RAM[7](44556677)/////////////
	///////////////////////////////////////////////
	///////////////////1_byte//////////////////////
	#1000 RX = 0;	      //開始02
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////2_byte//////////////////////
	#1000 RX = 0;       //開始 87(寫入ram[7])
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////3_byte//////////////////////
	#1000 RX = 0;       //開始 0100_0100
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////4_byte//////////////////////
	#1000 RX = 0;       //開始 0101_0101
	#1000 RX = 1;       
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////5_byte//////////////////////
	#1000 RX = 0;       //開始 0110_0110
	#1000 RX = 0;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////6_byte//////////////////////
	#1000 RX = 0;       //開始 0111_0111
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////7_byte//////////////////////
	#1000 RX = 0;       //開始 1100_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////8_byte//////////////////////
	#1000 RX = 0;       //開始 0000_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	#3000 RX = 1;
	///////////////////////////////////////////////
	////////////WRITE RAM[8](55667788)/////////////
	///////////////////////////////////////////////
	///////////////////1_byte//////////////////////
	#1000 RX = 0;	      //開始02
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////2_byte//////////////////////
	#1000 RX = 0;       //開始 88(寫入ram[8])
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////3_byte//////////////////////
	#1000 RX = 0;       //開始 0101_0101
	#1000 RX = 1;       
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////4_byte//////////////////////
	#1000 RX = 0;       //開始 0110_0110
	#1000 RX = 0;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////5_byte//////////////////////
	#1000 RX = 0;       //開始 0111_0111
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////6_byte//////////////////////
	#1000 RX = 0;       //開始 1000_1000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////7_byte//////////////////////
	#1000 RX = 0;       //開始 1100_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////8_byte//////////////////////
	#1000 RX = 0;       //開始 0000_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	#3000 RX = 1;
	///////////////////////////////
	//未寫完正確user_key時測試加密//
	///////////////////////////////
	///////////////////////////////////////////////
	////////////WRITE RAM[9](XXXXXXXX)/////////////
	///////////////////////////////////////////////
	///////////////////1_byte//////////////////////
	#1000 RX = 0;	      //開始02
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////2_byte//////////////////////
	#1000 RX = 0;       //開始 89(寫入ram[9])
	#1000 RX = 1;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////3_byte//////////////////////
	#1000 RX = 0;       //開始 0101_0101
	#1000 RX = 1;       
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////4_byte//////////////////////
	#1000 RX = 0;       //開始 0110_0110
	#1000 RX = 0;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////5_byte//////////////////////
	#1000 RX = 0;       //開始 0111_0111
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////6_byte//////////////////////
	#1000 RX = 0;       //開始 1000_1000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////7_byte//////////////////////
	#1000 RX = 0;       //開始 1100_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////8_byte//////////////////////
	#1000 RX = 0;       //開始 0000_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	#3000 RX = 1;
	////////////////////////////
	//寫完正確user_key後測試加密//
	////////////////////////////
	///////////////////////////////////////////////
	////////////WRITE RAM[24](F0DDCEDB)/////////////
	///////////////////////////////////////////////
	///////////////////1_byte//////////////////////
	#1000 RX = 0;	      //開始02
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////2_byte//////////////////////
	#1000 RX = 0;       //開始 98(寫入ram[24])
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////3_byte//////////////////////
	#1000 RX = 0;       //開始 1111_0000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////4_byte//////////////////////
	#1000 RX = 0;       //開始 1101_1101
	#1000 RX = 1;       
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////5_byte//////////////////////
	#1000 RX = 0;       //開始 1100_1110
	#1000 RX = 0;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////6_byte//////////////////////
	#1000 RX = 0;       //開始 1101_1011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////7_byte//////////////////////
	#1000 RX = 0;       //開始 1100_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////8_byte//////////////////////
	#1000 RX = 0;       //開始 0000_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	#3000 RX = 1;
	///////////////////////////////////////////////
	////////////WRITE RAM[9](XXXXXXXX)/////////////
	///////////////////////////////////////////////
	///////////////////1_byte//////////////////////
	#1000 RX = 0;	      //開始02
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////2_byte//////////////////////
	#1000 RX = 0;       //開始 89(寫入ram[9])
	#1000 RX = 1;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////3_byte//////////////////////
	#1000 RX = 0;       //開始 0101_0101
	#1000 RX = 1;       
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////4_byte//////////////////////
	#1000 RX = 0;       //開始 0110_0110
	#1000 RX = 0;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////5_byte//////////////////////
	#1000 RX = 0;       //開始 0111_0111
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////6_byte//////////////////////
	#1000 RX = 0;       //開始 1000_1000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////7_byte//////////////////////
	#1000 RX = 0;       //開始 1100_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////8_byte//////////////////////
	#1000 RX = 0;       //開始 0000_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	#3000 RX = 1;
	////////////////////////////
	//拿前面加密資料進行解密測試//
	////////////////////////////
	////////////////////////////
	///////////////////////////////////////////////
	////////////WRITE RAM[4](b0fdcae6)/////////////
	///////////////////////////////////////////////
	///////////////////1_byte//////////////////////
	#1000 RX = 0;	      //開始02
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////2_byte//////////////////////
	#1000 RX = 0;       //開始 84(寫入ram[4])
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////3_byte//////////////////////
	#1000 RX = 0;       //開始 b0 1011 0000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////4_byte//////////////////////
	#1000 RX = 0;       //開始 fd 1111 1101
	#1000 RX = 1;       
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////5_byte//////////////////////
	#1000 RX = 0;       //開始 ca 1100 1010
	#1000 RX = 0;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////6_byte//////////////////////
	#1000 RX = 0;       //開始 e6 1110 0110
	#1000 RX = 0;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////7_byte//////////////////////
	#1000 RX = 0;       //開始 1100_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////8_byte//////////////////////
	#1000 RX = 0;       //開始 0000_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	#3000 RX = 1;
	///////////////////////////////////////////////
	////////////WRITE RAM[5](8987d5b9)/////////////
	///////////////////////////////////////////////
	///////////////////1_byte//////////////////////
	#1000 RX = 0;	      //開始02
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////2_byte//////////////////////
	#1000 RX = 0;       //開始 85(寫入ram[5])
	#1000 RX = 1;       
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////3_byte//////////////////////
	#1000 RX = 0;       //開始 89 1000 1001
	#1000 RX = 1;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////4_byte//////////////////////
	#1000 RX = 0;       //開始 87 1000 0111
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////5_byte//////////////////////
	#1000 RX = 0;       //開始 d5 1101 0101
	#1000 RX = 1;       
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////6_byte//////////////////////
	#1000 RX = 0;       //開始 b9 1011 1001
	#1000 RX = 1;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////7_byte//////////////////////
	#1000 RX = 0;       //開始 1100_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////8_byte//////////////////////
	#1000 RX = 0;       //開始 0000_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	#3000 RX = 1;
	///////////////////////////////////////////////
	////////////WRITE RAM[6](e0a1dfc4)/////////////
	///////////////////////////////////////////////
	///////////////////1_byte//////////////////////
	#1000 RX = 0;	      //開始02
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////2_byte//////////////////////
	#1000 RX = 0;       //開始 86(寫入ram[6])
	#1000 RX = 0;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////3_byte//////////////////////
	#1000 RX = 0;       //開始 e0 1110 0000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////4_byte//////////////////////
	#1000 RX = 0;       //開始 a1 1010 0001
	#1000 RX = 1;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////5_byte//////////////////////
	#1000 RX = 0;       //開始 df 1101 1111
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////6_byte//////////////////////
	#1000 RX = 0;       //開始 c4 1100 0100
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////7_byte//////////////////////
	#1000 RX = 0;       //開始 1100_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////8_byte//////////////////////
	#1000 RX = 0;       //開始 0000_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	#3000 RX = 1;
	///////////////////////////////////////////////
	////////////WRITE RAM[7](8ea5ebe7)/////////////
	///////////////////////////////////////////////
	///////////////////1_byte//////////////////////
	#1000 RX = 0;	      //開始02
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////2_byte//////////////////////
	#1000 RX = 0;       //開始 87(寫入ram[7])
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////3_byte//////////////////////
	#1000 RX = 0;       //開始 8e 1000 1110
	#1000 RX = 0;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////4_byte//////////////////////
	#1000 RX = 0;       //開始 a5 1010 0101
	#1000 RX = 1;       
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////5_byte//////////////////////
	#1000 RX = 0;       //開始 eb 1110 1011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////6_byte//////////////////////
	#1000 RX = 0;       //開始 e7 1110 0111
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////7_byte//////////////////////
	#1000 RX = 0;       //開始 1100_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////8_byte//////////////////////
	#1000 RX = 0;       //開始 0000_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	#3000 RX = 1;
	///////////////////////////////////////////////
	////////////WRITE RAM[8](96c8feff)/////////////
	///////////////////////////////////////////////
	///////////////////1_byte//////////////////////
	#1000 RX = 0;	      //開始02
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////2_byte//////////////////////
	#1000 RX = 0;       //開始 88(寫入ram[8])
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////3_byte//////////////////////
	#1000 RX = 0;       //開始 96 1001 0110
	#1000 RX = 0;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////4_byte//////////////////////
	#1000 RX = 0;       //開始 c8 1100 1000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////5_byte//////////////////////
	#1000 RX = 0;       //開始 fe 1111 1110
	#1000 RX = 0;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////6_byte//////////////////////
	#1000 RX = 0;       //開始 ff
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////7_byte//////////////////////
	#1000 RX = 0;       //開始 1100_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////8_byte//////////////////////
	#1000 RX = 0;       //開始 0000_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	#3000 RX = 1;
	//////////////////////////////
	//未寫入正確user_key後測試解密//
	//////////////////////////////
	////////////////////////////////////////////////
	////////////WRITE RAM[24](00000000)/////////////
	///////////////////////////////////////////////
	///////////////////1_byte//////////////////////
	#1000 RX = 0;	      //開始02
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////2_byte//////////////////////
	#1000 RX = 0;       //開始 98(寫入ram[24])
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////3_byte//////////////////////
	#1000 RX = 0;       //開始 1000_0000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////4_byte//////////////////////
	#1000 RX = 0;       //開始 1000_0000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////5_byte//////////////////////
	#1000 RX = 0;       //開始 1000_0000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////6_byte//////////////////////
	#1000 RX = 0;       //開始 1000_0000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////7_byte//////////////////////
	#1000 RX = 0;       //開始 1100_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////8_byte//////////////////////
	#1000 RX = 0;       //開始 0000_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	#3000 RX = 1;
	///////////////////////////////////////////////
	////////////WRITE RAM[10](XXXXXXXX)/////////////
	///////////////////////////////////////////////
	///////////////////1_byte//////////////////////
	#1000 RX = 0;	      //開始02
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////2_byte//////////////////////
	#1000 RX = 0;       //開始 8a(寫入ram[10])
	#1000 RX = 0;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////3_byte//////////////////////
	#1000 RX = 0;       //開始 0101_0101
	#1000 RX = 1;       
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////4_byte//////////////////////
	#1000 RX = 0;       //開始 0110_0110
	#1000 RX = 0;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////5_byte//////////////////////
	#1000 RX = 0;       //開始 0111_0111
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////6_byte//////////////////////
	#1000 RX = 0;       //開始 1000_1000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////7_byte//////////////////////
	#1000 RX = 0;       //開始 1100_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////8_byte//////////////////////
	#1000 RX = 0;       //開始 0000_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	#6000 RX = 1;
	
	/////////////////////////////
	//寫入正確user_key後測試解密//
	/////////////////////////////
	/////////////////////////////
	///////////////////////////////////////////////
	////////////WRITE RAM[24](F0DDCEDB)/////////////
	///////////////////////////////////////////////
	///////////////////1_byte//////////////////////
	#1000 RX = 0;	      //開始02
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////2_byte//////////////////////
	#1000 RX = 0;       //開始 98(寫入ram[24])
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////3_byte//////////////////////
	#1000 RX = 0;       //開始 1111_0000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////4_byte//////////////////////
	#1000 RX = 0;       //開始 1101_1101
	#1000 RX = 1;       
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////5_byte//////////////////////
	#1000 RX = 0;       //開始 1100_1110
	#1000 RX = 0;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////6_byte//////////////////////
	#1000 RX = 0;       //開始 1101_1011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////7_byte//////////////////////
	#1000 RX = 0;       //開始 1100_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////8_byte//////////////////////
	#1000 RX = 0;       //開始 0000_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	#3000 RX = 1;
	///////////////////////////////////////////////
	////////////WRITE RAM[10](XXXXXXXX)/////////////
	///////////////////////////////////////////////
	///////////////////1_byte//////////////////////
	#1000 RX = 0;	      //開始02
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////2_byte//////////////////////
	#1000 RX = 0;       //開始 8a(寫入ram[10])
	#1000 RX = 0;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////3_byte//////////////////////
	#1000 RX = 0;       //開始 0101_0101
	#1000 RX = 1;       
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////4_byte//////////////////////
	#1000 RX = 0;       //開始 0110_0110
	#1000 RX = 0;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////5_byte//////////////////////
	#1000 RX = 0;       //開始 0111_0111
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////6_byte//////////////////////
	#1000 RX = 0;       //開始 1000_1000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////7_byte//////////////////////
	#1000 RX = 0;       //開始 1100_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////8_byte//////////////////////
	#1000 RX = 0;       //開始 0000_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	#20000 RX = 1;
	
	////////////
	////256/////
	////////////
	///////////////////////////////////////////////
	////////////WRITE RAM[29](80808081)/////////////
	///////////////////////////////////////////////
	///////////////////1_byte//////////////////////
	#1000 RX = 0;	      //開始02
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////2_byte//////////////////////
	#1000 RX = 0;       //開始 9D(寫入ram[29])
	#1000 RX = 1;       
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////3_byte//////////////////////
	#1000 RX = 0;       //開始 1000_0001
	#1000 RX = 1;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////4_byte//////////////////////
	#1000 RX = 0;       //開始 1000_0000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////5_byte//////////////////////
	#1000 RX = 0;       //開始 1000_0000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////6_byte//////////////////////
	#1000 RX = 0;       //開始 1000_0000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////7_byte//////////////////////
	#1000 RX = 0;       //開始 1100_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////8_byte//////////////////////
	#1000 RX = 0;       //開始 0000_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	#3000 RX = 1;
	///////////////////////////////////////////////
	////////////WRITE RAM[30](80808080)/////////////
	///////////////////////////////////////////////
	///////////////////1_byte//////////////////////
	#1000 RX = 0;	      //開始02
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////2_byte//////////////////////
	#1000 RX = 0;       //開始 9E(寫入ram[30])
	#1000 RX = 0;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////3_byte//////////////////////
	#1000 RX = 0;       //開始 1000_0000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////4_byte//////////////////////
	#1000 RX = 0;       //開始 1000_0000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////5_byte//////////////////////
	#1000 RX = 0;       //開始 1000_0000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////6_byte//////////////////////
	#1000 RX = 0;       //開始 1000_0000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////7_byte//////////////////////
	#1000 RX = 0;       //開始 1100_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////8_byte//////////////////////
	#1000 RX = 0;       //開始 0000_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	#3000 RX = 1;
	///////////////////////////////////////////////
	////////////WRITE RAM[31](80808080)/////////////
	///////////////////////////////////////////////
	///////////////////1_byte//////////////////////
	#1000 RX = 0;	      //開始02
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////2_byte//////////////////////
	#1000 RX = 0;       //開始 9F(寫入ram[31])
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////3_byte//////////////////////
	#1000 RX = 0;       //開始 1000_0000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////4_byte//////////////////////
	#1000 RX = 0;       //開始 1000_0000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////5_byte//////////////////////
	#1000 RX = 0;       //開始 1000_0000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////6_byte//////////////////////
	#1000 RX = 0;       //開始 1000_0000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////7_byte//////////////////////
	#1000 RX = 0;       //開始 1100_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////8_byte//////////////////////
	#1000 RX = 0;       //開始 0000_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	#3000 RX = 1;
	///////////////////////////////////////////////
	////////////WRITE RAM[32](80808080)/////////////
	///////////////////////////////////////////////
	///////////////////1_byte//////////////////////
	#1000 RX = 0;	      //開始02
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////2_byte//////////////////////
	#1000 RX = 0;       //開始 A0(寫入ram[32])
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////3_byte//////////////////////
	#1000 RX = 0;       //開始 1000_0000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////4_byte//////////////////////
	#1000 RX = 0;       //開始 1000_0000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////5_byte//////////////////////
	#1000 RX = 0;       //開始 1000_0000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////6_byte//////////////////////
	#1000 RX = 0;       //開始 1000_0000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////7_byte//////////////////////
	#1000 RX = 0;       //開始 1100_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////8_byte//////////////////////
	#1000 RX = 0;       //開始 0000_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	#3000 RX = 1;
	///////////////////////////////////////////////
	////////////WRITE RAM[33](81808080)/////////////
	///////////////////////////////////////////////
	///////////////////1_byte//////////////////////
	#1000 RX = 0;	      //開始02
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////2_byte//////////////////////
	#1000 RX = 0;       //開始 A1(寫入ram[33])
	#1000 RX = 1;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////3_byte//////////////////////
	#1000 RX = 0;       //開始 1000_0001
	#1000 RX = 1;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////4_byte//////////////////////
	#1000 RX = 0;       //開始 1000_0000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////5_byte//////////////////////
	#1000 RX = 0;       //開始 1000_0000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////6_byte//////////////////////
	#1000 RX = 0;       //開始 1000_0000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////7_byte//////////////////////
	#1000 RX = 0;       //開始 1100_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////8_byte//////////////////////
	#1000 RX = 0;       //開始 0000_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	#3000 RX = 1;
	///////////////////////////
	/////未寫正確256key加密/////
	///////////////////////////////////////////////
	////////////WRITE RAM[11](XXXXXXXX)/////////////
	///////////////////////////////////////////////
	///////////////////1_byte//////////////////////
	#1000 RX = 0;	      //開始02
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////2_byte//////////////////////
	#1000 RX = 0;       //開始 8b(寫入ram[11])
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////3_byte//////////////////////
	#1000 RX = 0;       //開始 0101_0101
	#1000 RX = 1;       
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////4_byte//////////////////////
	#1000 RX = 0;       //開始 0110_0110
	#1000 RX = 0;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////5_byte//////////////////////
	#1000 RX = 0;       //開始 0111_0111
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////6_byte//////////////////////
	#1000 RX = 0;       //開始 1000_1000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////7_byte//////////////////////
	#1000 RX = 0;       //開始 1100_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////8_byte//////////////////////
	#1000 RX = 0;       //開始 0000_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	#3000 RX = 1;
	///////////////////////////////////////////////
	////////////WRITE RAM[33](80808080)/////////////
	///////////////////////////////////////////////
	///////////////////1_byte//////////////////////
	#1000 RX = 0;	      //開始02
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////2_byte//////////////////////
	#1000 RX = 0;       //開始 A1(寫入ram[33])
	#1000 RX = 1;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////3_byte//////////////////////
	#1000 RX = 0;       //開始 1000_0000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////4_byte//////////////////////
	#1000 RX = 0;       //開始 1000_0000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////5_byte//////////////////////
	#1000 RX = 0;       //開始 1000_0000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////6_byte//////////////////////
	#1000 RX = 0;       //開始 1000_0000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////7_byte//////////////////////
	#1000 RX = 0;       //開始 1100_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////8_byte//////////////////////
	#1000 RX = 0;       //開始 0000_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	#3000 RX = 1;
	////////////////////////////
	/////寫正確256key加密/////////
	///////////////////////////////////////////////
	////////////WRITE RAM[11](XXXXXXXX)/////////////
	///////////////////////////////////////////////
	///////////////////1_byte//////////////////////
	#1000 RX = 0;	      //開始02
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////2_byte//////////////////////
	#1000 RX = 0;       //開始 8b(寫入ram[11])
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////3_byte//////////////////////
	#1000 RX = 0;       //開始 0101_0101
	#1000 RX = 1;       
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////4_byte//////////////////////
	#1000 RX = 0;       //開始 0110_0110
	#1000 RX = 0;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////5_byte//////////////////////
	#1000 RX = 0;       //開始 0111_0111
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////6_byte//////////////////////
	#1000 RX = 0;       //開始 1000_1000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////7_byte//////////////////////
	#1000 RX = 0;       //開始 1100_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////8_byte//////////////////////
	#1000 RX = 0;       //開始 0000_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	#20000 RX = 1;
	
	
	////////////////////////////
	//拿前面加密資料進行解密測試//
	////////////////////////////
	////////////////////////////
	///////////////////////////////////////////////
	////////////WRITE RAM[4](b3e8c5ee)/////////////
	///////////////////////////////////////////////
	///////////////////1_byte//////////////////////
	#1000 RX = 0;	      //開始02
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////2_byte//////////////////////
	#1000 RX = 0;       //開始 84(寫入ram[4])
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////3_byte//////////////////////
	#1000 RX = 0;       //開始 b3 1011 0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////4_byte//////////////////////
	#1000 RX = 0;       //開始 e8 1110 1000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////5_byte//////////////////////
	#1000 RX = 0;       //開始 c5 1100 0101
	#1000 RX = 1;       
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////6_byte//////////////////////
	#1000 RX = 0;       //開始 ee 1110 1110
	#1000 RX = 0;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////7_byte//////////////////////
	#1000 RX = 0;       //開始 1100_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////8_byte//////////////////////
	#1000 RX = 0;       //開始 0000_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	#3000 RX = 1;
	///////////////////////////////////////////////
	////////////WRITE RAM[5](caf6e5b8)/////////////
	///////////////////////////////////////////////
	///////////////////1_byte//////////////////////
	#1000 RX = 0;	      //開始02
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////2_byte//////////////////////
	#1000 RX = 0;       //開始 85(寫入ram[5])
	#1000 RX = 1;       
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////3_byte//////////////////////
	#1000 RX = 0;       //開始 ca 1100 1010
	#1000 RX = 0;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////4_byte//////////////////////
	#1000 RX = 0;       //開始 f6 1111 0110
	#1000 RX = 0;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////5_byte//////////////////////
	#1000 RX = 0;       //開始  e5 1110 0101
	#1000 RX = 1;       
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////6_byte//////////////////////
	#1000 RX = 0;       //開始 b8 1011 1000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////7_byte//////////////////////
	#1000 RX = 0;       //開始 1100_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////8_byte//////////////////////
	#1000 RX = 0;       //開始 0000_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	#3000 RX = 1;
	///////////////////////////////////////////////
	////////////WRITE RAM[6](978ce992)/////////////
	///////////////////////////////////////////////
	///////////////////1_byte//////////////////////
	#1000 RX = 0;	      //開始02
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////2_byte//////////////////////
	#1000 RX = 0;       //開始 86(寫入ram[6])
	#1000 RX = 0;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////3_byte//////////////////////
	#1000 RX = 0;       //開始 97 1001 0111
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////4_byte//////////////////////
	#1000 RX = 0;       //開始 8c 1000 1100
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////5_byte//////////////////////
	#1000 RX = 0;       //開始 e9 1110 1001
	#1000 RX = 1;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////6_byte//////////////////////
	#1000 RX = 0;       //開始 92 1001 0010
	#1000 RX = 0;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////7_byte//////////////////////
	#1000 RX = 0;       //開始 1100_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////8_byte//////////////////////
	#1000 RX = 0;       //開始 0000_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	#3000 RX = 1;
	///////////////////////////////////////////////
	////////////WRITE RAM[7](b3adf290)/////////////
	///////////////////////////////////////////////
	///////////////////1_byte//////////////////////
	#1000 RX = 0;	      //開始02
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////2_byte//////////////////////
	#1000 RX = 0;       //開始 87(寫入ram[7])
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////3_byte//////////////////////
	#1000 RX = 0;       //開始 b3 1011 0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////4_byte//////////////////////
	#1000 RX = 0;       //開始 ad 1010 1101
	#1000 RX = 1;       
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////5_byte//////////////////////
	#1000 RX = 0;       //開始 f2 1111 0010
	#1000 RX = 0;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////6_byte//////////////////////
	#1000 RX = 0;       //開始 90 1001 0000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////7_byte//////////////////////
	#1000 RX = 0;       //開始 1100_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////8_byte//////////////////////
	#1000 RX = 0;       //開始 0000_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	#3000 RX = 1;
	///////////////////////////////////////////////
	////////////WRITE RAM[8](db80fcff)/////////////
	///////////////////////////////////////////////
	///////////////////1_byte//////////////////////
	#1000 RX = 0;	      //開始02
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////2_byte//////////////////////
	#1000 RX = 0;       //開始 88(寫入ram[8])
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////3_byte//////////////////////
	#1000 RX = 0;       //開始 db 1101 1011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////4_byte//////////////////////
	#1000 RX = 0;       //開始 80 1000 0000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////5_byte//////////////////////
	#1000 RX = 0;       //開始 fc 1111 1100
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////6_byte//////////////////////
	#1000 RX = 0;       //開始 ff 1111 1111
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////7_byte//////////////////////
	#1000 RX = 0;       //開始 1100_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////8_byte//////////////////////
	#1000 RX = 0;       //開始 0000_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	#3000 RX = 1;
	//////////////////////////////
	//未寫入正確user_key後測試解密//
	//////////////////////////////
	////////////////////////////////////////////////
	////////////WRITE RAM[24](00000000)/////////////
	///////////////////////////////////////////////
	///////////////////1_byte//////////////////////
	#1000 RX = 0;	      //開始02
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////2_byte//////////////////////
	#1000 RX = 0;       //開始 98(寫入ram[24])
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////3_byte//////////////////////
	#1000 RX = 0;       //開始 1000_0000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////4_byte//////////////////////
	#1000 RX = 0;       //開始 1000_0000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////5_byte//////////////////////
	#1000 RX = 0;       //開始 1000_0000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////6_byte//////////////////////
	#1000 RX = 0;       //開始 1000_0000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////7_byte//////////////////////
	#1000 RX = 0;       //開始 1100_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////8_byte//////////////////////
	#1000 RX = 0;       //開始 0000_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	#3000 RX = 1;
	///////////////////////////////////////////////
	////////////WRITE RAM[12](XXXXXXXX)/////////////
	///////////////////////////////////////////////
	///////////////////1_byte//////////////////////
	#1000 RX = 0;	      //開始02
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////2_byte//////////////////////
	#1000 RX = 0;       //開始 8c(寫入ram[12])
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////3_byte//////////////////////
	#1000 RX = 0;       //開始 0101_0101
	#1000 RX = 1;       
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////4_byte//////////////////////
	#1000 RX = 0;       //開始 0110_0110
	#1000 RX = 0;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////5_byte//////////////////////
	#1000 RX = 0;       //開始 0111_0111
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////6_byte//////////////////////
	#1000 RX = 0;       //開始 1000_1000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////7_byte//////////////////////
	#1000 RX = 0;       //開始 1100_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////8_byte//////////////////////
	#1000 RX = 0;       //開始 0000_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	#6000 RX = 1;
	
	/////////////////////////////
	//寫入正確user_key後測試解密//
	/////////////////////////////
	/////////////////////////////
	///////////////////////////////////////////////
	////////////WRITE RAM[24](F0DDCEDB)/////////////
	///////////////////////////////////////////////
	///////////////////1_byte//////////////////////
	#1000 RX = 0;	      //開始02
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////2_byte//////////////////////
	#1000 RX = 0;       //開始 98(寫入ram[24])
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////3_byte//////////////////////
	#1000 RX = 0;       //開始 1111_0000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////4_byte//////////////////////
	#1000 RX = 0;       //開始 1101_1101
	#1000 RX = 1;       
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////5_byte//////////////////////
	#1000 RX = 0;       //開始 1100_1110
	#1000 RX = 0;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////6_byte//////////////////////
	#1000 RX = 0;       //開始 1101_1011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////7_byte//////////////////////
	#1000 RX = 0;       //開始 1100_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////8_byte//////////////////////
	#1000 RX = 0;       //開始 0000_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	#3000 RX = 1;
	///////////////////////////////////////////////
	////////////WRITE RAM[12](XXXXXXXX)/////////////
	///////////////////////////////////////////////
	///////////////////1_byte//////////////////////
	#1000 RX = 0;	      //開始02
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////2_byte//////////////////////
	#1000 RX = 0;       //開始 8c(寫入ram[12])
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////3_byte//////////////////////
	#1000 RX = 0;       //開始 0101_0101
	#1000 RX = 1;       
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////4_byte//////////////////////
	#1000 RX = 0;       //開始 0110_0110
	#1000 RX = 0;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////5_byte//////////////////////
	#1000 RX = 0;       //開始 0111_0111
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////6_byte//////////////////////
	#1000 RX = 0;       //開始 1000_1000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////7_byte//////////////////////
	#1000 RX = 0;       //開始 1100_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////8_byte//////////////////////
	#1000 RX = 0;       //開始 0000_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	#800000 RX = 1;
	
	////////////////////////////////////////////////
	
	#250000 $stop;      //執行到指定時間後停止
	end
  
	always #10 clk = ~clk;
  
endmodule



