library verilog;
use verilog.vl_types.all;
entity AES_tb is
end AES_tb;
