library verilog;
use verilog.vl_types.all;
entity rs232_test is
end rs232_test;
