library verilog;
use verilog.vl_types.all;
entity inverseMixColumns is
    port(
        state_in        : in     vl_logic_vector(127 downto 0);
        state_out       : out    vl_logic_vector(127 downto 0)
    );
end inverseMixColumns;
