module bits64_test;
  
	wire TX;
	reg  RX, clk, rst, sw2, sw1 ,sw0;
	wire [7:0]port_b_out;
  
	rs232 f_rs232(TX, RX, sw2, sw1 ,sw0, clk, rst, port_b_out);
	initial begin
		rst = 1; clk = 0; RX = 1; sw2 = 0; sw1 = 0; sw0 = 0; //按下reset並將clk清0
	#20 rst = 0;  		   //放開reset
  ///////////////////////////////////////////////
  ///////////////////測試非02開始/////////////////
  ///////////////////////////////////////////////
  
	#890 RX = 0;	      //開始0100_0000
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 1;
	#890 RX = 0;
	#890 RX = 1;       //結束(非02因此未開始)
	#3000 RX = 1;
	
	///////////////////////////////////////////////
  ///////////////測試8bytes但非03結束/////////////
  ///////////////////////////////////////////////
  
	///////////////////1_byte//////////////////////
	#890 RX = 0;	      //開始0000_0010
	#890 RX = 0;
	#890 RX = 1;
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 1;       //結束
	///////////////////2_byte//////////////////////
	#890 RX = 0;       //開始 1111_1111
	#890 RX = 1;       
	#890 RX = 1;
	#890 RX = 1;
	#890 RX = 1;
	#890 RX = 1;
	#890 RX = 1;
	#890 RX = 1;
	#890 RX = 1;
	#890 RX = 1;       //結束
	///////////////////3_byte//////////////////////
	#890 RX = 0;       //開始 1111_0000
	#890 RX = 0;       
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 1;
	#890 RX = 1;
	#890 RX = 1;
	#890 RX = 1;
	#890 RX = 1;       //結束
	///////////////////4_byte//////////////////////
	#890 RX = 0;       //開始 0101_0101
	#890 RX = 1;       
	#890 RX = 0;
	#890 RX = 1;
	#890 RX = 0;
	#890 RX = 1;
	#890 RX = 0;
	#890 RX = 1;
	#890 RX = 0;
	#890 RX = 1;       //結束
	///////////////////5_byte//////////////////////
	#890 RX = 0;       //開始 1010_1010
	#890 RX = 0;       
	#890 RX = 1;
	#890 RX = 0;
	#890 RX = 1;
	#890 RX = 0;
	#890 RX = 1;
	#890 RX = 0;
	#890 RX = 1;
	#890 RX = 1;       //結束
	///////////////////6_byte//////////////////////
	#890 RX = 0;       //開始 0011_1100
	#890 RX = 0;       
	#890 RX = 0;
	#890 RX = 1;
	#890 RX = 1;
	#890 RX = 1;
	#890 RX = 1;
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 1;       //結束
	///////////////////7_byte//////////////////////
	#890 RX = 0;       //開始 1100_0011
	#890 RX = 1;       
	#890 RX = 1;
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 1;
	#890 RX = 1;
	#890 RX = 1;       //結束
	///////////////////8_byte//////////////////////
	#890 RX = 0;       //開始 1100_0000
	#890 RX = 0;       
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 1;
	#890 RX = 1;
	#890 RX = 1;       //結束
	#5000 RX = 1;
	
	
	///////////////////////////////////////////////
  //////////////測試正確8bytes(寫入)//////////////
  ///////////////////////////////////////////////
	
	///////////////////1_byte//////////////////////
	#890 RX = 0;	      //開始0000_0010
	#890 RX = 0;
	#890 RX = 1;
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 1;       //結束
	///////////////////2_byte//////////////////////
	#890 RX = 0;       //開始 1111_1111
	#890 RX = 1;       
	#890 RX = 1;
	#890 RX = 1;
	#890 RX = 1;
	#890 RX = 1;
	#890 RX = 1;
	#890 RX = 1;
	#890 RX = 1;
	#890 RX = 1;       //結束
	///////////////////3_byte//////////////////////
	#890 RX = 0;       //開始 1111_0000
	#890 RX = 0;       
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 1;
	#890 RX = 1;
	#890 RX = 1;
	#890 RX = 1;
	#890 RX = 1;       //結束
	///////////////////4_byte//////////////////////
	#890 RX = 0;       //開始 0101_0101
	#890 RX = 1;       
	#890 RX = 0;
	#890 RX = 1;
	#890 RX = 0;
	#890 RX = 1;
	#890 RX = 0;
	#890 RX = 1;
	#890 RX = 0;
	#890 RX = 1;       //結束
	///////////////////5_byte//////////////////////
	#890 RX = 0;       //開始 1010_1010
	#890 RX = 0;       
	#890 RX = 1;
	#890 RX = 0;
	#890 RX = 1;
	#890 RX = 0;
	#890 RX = 1;
	#890 RX = 0;
	#890 RX = 1;
	#890 RX = 1;       //結束
	///////////////////6_byte//////////////////////
	#890 RX = 0;       //開始 0011_1100
	#890 RX = 0;       
	#890 RX = 0;
	#890 RX = 1;
	#890 RX = 1;
	#890 RX = 1;
	#890 RX = 1;
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 1;       //結束
	///////////////////7_byte//////////////////////
	#890 RX = 0;       //開始 1100_0011
	#890 RX = 1;       
	#890 RX = 1;
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 1;
	#890 RX = 1;
	#890 RX = 1;       //結束
	///////////////////8_byte//////////////////////
	#890 RX = 0;       //開始 0000_0011
	#890 RX = 1;       
	#890 RX = 1;
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 1;       //結束
	#3000 RX = 1;
	
	///////////////////////////////////////////////
  //////////////寫(掉)//////////////
  ///////////////////////////////////////////////
	
	///////////////////1_byte//////////////////////
	#890 RX = 0;	      //開始0000_0010
	#890 RX = 0;
	#890 RX = 1;
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 1;       //結束
	///////////////////2_byte//////////////////////
	#890 RX = 0;       //開始 1111_1111
	#890 RX = 1;       
	#890 RX = 1;
	#890 RX = 1;
	#890 RX = 1;
	#890 RX = 1;
	#890 RX = 1;
	#890 RX = 1;
	#890 RX = 1;
	#890 RX = 1;       //結束
	///////////////////3_byte//////////////////////
	#890 RX = 0;       //開始 1111_0000
	#890 RX = 0;       
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 1;
	#890 RX = 1;
	#890 RX = 1;
	#890 RX = 1;
	#890 RX = 1;       //結束
	///////////////////4_byte//////////////////////
	#890 RX = 0;       //開始 0101_0101
	#890 RX = 1;       
	#890 RX = 0;
	#890 RX = 1;
	#890 RX = 0;
	#890 RX = 1;
	#890 RX = 0;
	#890 RX = 1;
	#890 RX = 0;
	#890 RX = 1;       //結束
	///////////////////5_byte//////////////////////
	//掉
	///////////////////6_byte//////////////////////
	#890 RX = 0;       //開始 0011_1100
	#890 RX = 0;       
	#890 RX = 0;
	#890 RX = 1;
	#890 RX = 1;
	#890 RX = 1;
	#890 RX = 1;
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 1;       //結束
	///////////////////7_byte//////////////////////
	#890 RX = 0;       //開始 1100_0011
	#890 RX = 1;       
	#890 RX = 1;
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 1;
	#890 RX = 1;
	#890 RX = 1;       //結束
	///////////////////8_byte//////////////////////
	#890 RX = 0;       //開始 0000_1111
	#890 RX = 1;       
	#890 RX = 1;
	#890 RX = 1;
	#890 RX = 1;
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 1;       //結束
	#80000 RX = 1;
	
	#890 RX = 0;       //開始 0000_0011
	#890 RX = 1;       
	#890 RX = 1;
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 1;       //結束
	///////////////////////////////////////////////
  //////////////測試正確8bytes(讀取)//////////////
  ///////////////////////////////////////////////
	
	///////////////////1_byte//////////////////////
	#890 RX = 0;	      //開始0000_0010
	#890 RX = 0;
	#890 RX = 1;
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 1;       //結束
	///////////////////2_byte//////////////////////
	#890 RX = 0;       //開始 0111_1111
	#890 RX = 1;       
	#890 RX = 1;
	#890 RX = 1;
	#890 RX = 1;
	#890 RX = 1;
	#890 RX = 1;
	#890 RX = 1;
	#890 RX = 0;
	#890 RX = 1;       //結束
	///////////////////3_byte//////////////////////
	#890 RX = 0;       //開始 1111_0000
	#890 RX = 0;       
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 1;
	#890 RX = 1;
	#890 RX = 1;
	#890 RX = 1;
	#890 RX = 1;       //結束
	///////////////////4_byte//////////////////////
	#890 RX = 0;       //開始 0101_0101
	#890 RX = 1;       
	#890 RX = 0;
	#890 RX = 1;
	#890 RX = 0;
	#890 RX = 1;
	#890 RX = 0;
	#890 RX = 1;
	#890 RX = 0;
	#890 RX = 1;       //結束
	///////////////////5_byte//////////////////////
	#890 RX = 0;       //開始 1010_1010
	#890 RX = 0;       
	#890 RX = 1;
	#890 RX = 0;
	#890 RX = 1;
	#890 RX = 0;
	#890 RX = 1;
	#890 RX = 0;
	#890 RX = 1;
	#890 RX = 1;       //結束
	///////////////////6_byte//////////////////////
	#890 RX = 0;       //開始 0011_1100
	#890 RX = 0;       
	#890 RX = 0;
	#890 RX = 1;
	#890 RX = 1;
	#890 RX = 1;
	#890 RX = 1;
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 1;       //結束
	///////////////////7_byte//////////////////////
	#890 RX = 0;       //開始 1100_0011
	#890 RX = 1;       
	#890 RX = 1;
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 1;
	#890 RX = 1;
	#890 RX = 1;       //結束
	///////////////////8_byte//////////////////////
	#890 RX = 0;       //開始 0000_0011
	#890 RX = 1;       
	#890 RX = 1;
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 0;
	#890 RX = 1;       //結束
	
	#2000 sw2=0;sw1=0;sw0=1;
	#2000 sw2=0;sw1=1;sw0=0;
	#2000 sw2=0;sw1=1;sw0=1;
	///////////////////////////////////////////////////
	
	#80000 $stop;      //執行到指定時間後停止
	end
  
	always #10 clk = ~clk;
  
endmodule

