library verilog;
use verilog.vl_types.all;
entity bits64_test is
end bits64_test;
