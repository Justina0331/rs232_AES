module aes_data_tb;
  
	wire TX;
	reg  RX, clk, rst;
  
	rs232 f_rs232(TX, RX, clk, rst);
	initial begin
		rst = 1; clk = 0; RX = 1; //按下reset並將clk清0
	#20 rst = 0;  		   //放開reset
	
	///////////////////
	///////寫入DATA////
	///////////////////
	///////////////////////////////////////////////
	////////////WRITE RAM[4](11223344)/////////////
	///////////////////////////////////////////////
	///////////////////1_byte//////////////////////
	#1000 RX = 0;	      //開始02
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////2_byte//////////////////////
	#1000 RX = 0;       //開始 84(寫入ram[4])
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////3_byte//////////////////////
	#1000 RX = 0;       //開始 0001_0001
	#1000 RX = 1;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////4_byte//////////////////////
	#1000 RX = 0;       //開始 0010_0010
	#1000 RX = 0;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////5_byte//////////////////////
	#1000 RX = 0;       //開始 0011_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////6_byte//////////////////////
	#1000 RX = 0;       //開始 0100_0100
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////7_byte//////////////////////
	#1000 RX = 0;       //開始 1100_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////8_byte//////////////////////
	#1000 RX = 0;       //開始 0000_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	#3000 RX = 1;
	///////////////////////////////////////////////
	////////////WRITE RAM[5](22334455)/////////////
	///////////////////////////////////////////////
	///////////////////1_byte//////////////////////
	#1000 RX = 0;	      //開始02
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////2_byte//////////////////////
	#1000 RX = 0;       //開始 85(寫入ram[5])
	#1000 RX = 1;       
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////3_byte//////////////////////
	#1000 RX = 0;       //開始 0010_0010
	#1000 RX = 0;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////4_byte//////////////////////
	#1000 RX = 0;       //開始 0011_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////5_byte//////////////////////
	#1000 RX = 0;       //開始 0100_0100
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////6_byte//////////////////////
	#1000 RX = 0;       //開始 0101_0101
	#1000 RX = 1;       
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////7_byte//////////////////////
	#1000 RX = 0;       //開始 1100_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////8_byte//////////////////////
	#1000 RX = 0;       //開始 0000_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	#3000 RX = 1;
	///////////////////////////////////////////////
	////////////WRITE RAM[6](33445566)/////////////
	///////////////////////////////////////////////
	///////////////////1_byte//////////////////////
	#1000 RX = 0;	      //開始02
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////2_byte//////////////////////
	#1000 RX = 0;       //開始 86(寫入ram[6])
	#1000 RX = 0;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////3_byte//////////////////////
	#1000 RX = 0;       //開始 0011_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////4_byte//////////////////////
	#1000 RX = 0;       //開始 0100_0100
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////5_byte//////////////////////
	#1000 RX = 0;       //開始 0101_0101
	#1000 RX = 1;       
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////6_byte//////////////////////
	#1000 RX = 0;       //開始 0110_0110
	#1000 RX = 0;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////7_byte//////////////////////
	#1000 RX = 0;       //開始 1100_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////8_byte//////////////////////
	#1000 RX = 0;       //開始 0000_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	#3000 RX = 1;
	///////////////////////////////////////////////
	////////////WRITE RAM[7](44556677)/////////////
	///////////////////////////////////////////////
	///////////////////1_byte//////////////////////
	#1000 RX = 0;	      //開始02
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////2_byte//////////////////////
	#1000 RX = 0;       //開始 87(寫入ram[7])
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////3_byte//////////////////////
	#1000 RX = 0;       //開始 0100_0100
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////4_byte//////////////////////
	#1000 RX = 0;       //開始 0101_0101
	#1000 RX = 1;       
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////5_byte//////////////////////
	#1000 RX = 0;       //開始 0110_0110
	#1000 RX = 0;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////6_byte//////////////////////
	#1000 RX = 0;       //開始 0111_0111
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////7_byte//////////////////////
	#1000 RX = 0;       //開始 1100_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////8_byte//////////////////////
	#1000 RX = 0;       //開始 0000_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	#3000 RX = 1;
	///////////////////////////////////////////////
	////////////WRITE RAM[8](55667788)/////////////
	///////////////////////////////////////////////
	///////////////////1_byte//////////////////////
	#1000 RX = 0;	      //開始02
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////2_byte//////////////////////
	#1000 RX = 0;       //開始 88(寫入ram[8])
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////3_byte//////////////////////
	#1000 RX = 0;       //開始 0101_0101
	#1000 RX = 1;       
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////4_byte//////////////////////
	#1000 RX = 0;       //開始 0110_0110
	#1000 RX = 0;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////5_byte//////////////////////
	#1000 RX = 0;       //開始 0111_0111
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////6_byte//////////////////////
	#1000 RX = 0;       //開始 1000_1000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////7_byte//////////////////////
	#1000 RX = 0;       //開始 1100_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////8_byte//////////////////////
	#1000 RX = 0;       //開始 0000_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	#3000 RX = 1;
	///////////////////////////////////////////////
	////////////WRITE RAM[9](XXXXXXXX)/////////////
	///////////////////////////////////////////////
	///////////////////1_byte//////////////////////
	#1000 RX = 0;	      //開始02
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////2_byte//////////////////////
	#1000 RX = 0;       //開始 89(寫入ram[9])
	#1000 RX = 1;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////3_byte//////////////////////
	#1000 RX = 0;       //開始 0101_0101
	#1000 RX = 1;       
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////4_byte//////////////////////
	#1000 RX = 0;       //開始 0110_0110
	#1000 RX = 0;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////5_byte//////////////////////
	#1000 RX = 0;       //開始 0111_0111
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////6_byte//////////////////////
	#1000 RX = 0;       //開始 1000_1000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////7_byte//////////////////////
	#1000 RX = 0;       //開始 1100_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////8_byte//////////////////////
	#1000 RX = 0;       //開始 0000_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	#3000 RX = 1;
	
	
	
	////////////////////////////
	//拿前面加密資料進行解密測試//
	////////////////////////////
	//////////////////
	///////////////////////////////////////////////
	////////////WRITE RAM[4](b0fdcae6)/////////////
	///////////////////////////////////////////////
	///////////////////1_byte//////////////////////
	#1000 RX = 0;	      //開始02
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////2_byte//////////////////////
	#1000 RX = 0;       //開始 84(寫入ram[4])
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////3_byte//////////////////////
	#1000 RX = 0;       //開始 b0 1011 0000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////4_byte//////////////////////
	#1000 RX = 0;       //開始 fd 1111 1101
	#1000 RX = 1;       
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////5_byte//////////////////////
	#1000 RX = 0;       //開始 ca 1100 1010
	#1000 RX = 0;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////6_byte//////////////////////
	#1000 RX = 0;       //開始 e6 1110 0110
	#1000 RX = 0;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////7_byte//////////////////////
	#1000 RX = 0;       //開始 1100_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////8_byte//////////////////////
	#1000 RX = 0;       //開始 0000_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	#3000 RX = 1;
	///////////////////////////////////////////////
	////////////WRITE RAM[5](8987d5b9)/////////////
	///////////////////////////////////////////////
	///////////////////1_byte//////////////////////
	#1000 RX = 0;	      //開始02
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////2_byte//////////////////////
	#1000 RX = 0;       //開始 85(寫入ram[5])
	#1000 RX = 1;       
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////3_byte//////////////////////
	#1000 RX = 0;       //開始 89 1000 1001
	#1000 RX = 1;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////4_byte//////////////////////
	#1000 RX = 0;       //開始 87 1000 0111
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////5_byte//////////////////////
	#1000 RX = 0;       //開始 d5 1101 0101
	#1000 RX = 1;       
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////6_byte//////////////////////
	#1000 RX = 0;       //開始 b9 1011 1001
	#1000 RX = 1;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////7_byte//////////////////////
	#1000 RX = 0;       //開始 1100_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////8_byte//////////////////////
	#1000 RX = 0;       //開始 0000_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	#3000 RX = 1;
	///////////////////////////////////////////////
	////////////WRITE RAM[6](e0a1dfc4)/////////////
	///////////////////////////////////////////////
	///////////////////1_byte//////////////////////
	#1000 RX = 0;	      //開始02
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////2_byte//////////////////////
	#1000 RX = 0;       //開始 86(寫入ram[6])
	#1000 RX = 0;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////3_byte//////////////////////
	#1000 RX = 0;       //開始 e0 1110 0000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////4_byte//////////////////////
	#1000 RX = 0;       //開始 a1 1010 0001
	#1000 RX = 1;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////5_byte//////////////////////
	#1000 RX = 0;       //開始 df 1101 1111
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////6_byte//////////////////////
	#1000 RX = 0;       //開始 c4 1100 0100
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////7_byte//////////////////////
	#1000 RX = 0;       //開始 1100_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////8_byte//////////////////////
	#1000 RX = 0;       //開始 0000_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	#3000 RX = 1;
	///////////////////////////////////////////////
	////////////WRITE RAM[7](8ea5ebe7)/////////////
	///////////////////////////////////////////////
	///////////////////1_byte//////////////////////
	#1000 RX = 0;	      //開始02
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////2_byte//////////////////////
	#1000 RX = 0;       //開始 87(寫入ram[7])
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////3_byte//////////////////////
	#1000 RX = 0;       //開始 8e 1000 1110
	#1000 RX = 0;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////4_byte//////////////////////
	#1000 RX = 0;       //開始 a5 1010 0101
	#1000 RX = 1;       
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////5_byte//////////////////////
	#1000 RX = 0;       //開始 eb 1110 1011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////6_byte//////////////////////
	#1000 RX = 0;       //開始 e7 1110 0111
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////7_byte//////////////////////
	#1000 RX = 0;       //開始 1100_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////8_byte//////////////////////
	#1000 RX = 0;       //開始 0000_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	#3000 RX = 1;
	///////////////////////////////////////////////
	////////////WRITE RAM[8](96c8feff)/////////////
	///////////////////////////////////////////////
	///////////////////1_byte//////////////////////
	#1000 RX = 0;	      //開始02
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////2_byte//////////////////////
	#1000 RX = 0;       //開始 88(寫入ram[8])
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////3_byte//////////////////////
	#1000 RX = 0;       //開始 96 1001 0110
	#1000 RX = 0;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////4_byte//////////////////////
	#1000 RX = 0;       //開始 c8 1100 1000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////5_byte//////////////////////
	#1000 RX = 0;       //開始 fe 1111 1110
	#1000 RX = 0;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////6_byte//////////////////////
	#1000 RX = 0;       //開始 ff
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////7_byte//////////////////////
	#1000 RX = 0;       //開始 1100_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////8_byte//////////////////////
	#1000 RX = 0;       //開始 0000_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	#3000 RX = 1;
	///////////////////////////////////////////////
	////////////WRITE RAM[10](XXXXXXXX)/////////////
	///////////////////////////////////////////////
	///////////////////1_byte//////////////////////
	#1000 RX = 0;	      //開始02
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////2_byte//////////////////////
	#1000 RX = 0;       //開始 8a(寫入ram[10])
	#1000 RX = 0;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////3_byte//////////////////////
	#1000 RX = 0;       //開始 0101_0101
	#1000 RX = 1;       
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////4_byte//////////////////////
	#1000 RX = 0;       //開始 0110_0110
	#1000 RX = 0;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////5_byte//////////////////////
	#1000 RX = 0;       //開始 0111_0111
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////6_byte//////////////////////
	#1000 RX = 0;       //開始 1000_1000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////7_byte//////////////////////
	#1000 RX = 0;       //開始 1100_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////8_byte//////////////////////
	#1000 RX = 0;       //開始 0000_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	#60000 RX = 1;
	
	
	
	
	/*
	
	///////////////////////////////////////////////
	//////測試正確8bytes(讀出RAM[64](aes_RAM[1]))//////
	///////////////////////////////////////////////
	
	///////////////////1_byte//////////////////////
	#1000 RX = 0;	      //開始02
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////2_byte//////////////////////
	#1000 RX = 0;       //開始 40(讀出ram[64])0100 0000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////3_byte//////////////////////
	#1000 RX = 0;       //開始 0101_0101
	#1000 RX = 1;       
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////4_byte//////////////////////
	#1000 RX = 0;       //開始 0110_0110
	#1000 RX = 0;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////5_byte//////////////////////
	#1000 RX = 0;       //開始 0111_0111
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////6_byte//////////////////////
	#1000 RX = 0;       //開始 1000_1000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////7_byte//////////////////////
	#1000 RX = 0;       //開始 1100_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////8_byte//////////////////////
	#1000 RX = 0;       //開始 0000_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	#3000 RX = 1;
	
	////////////////////////////////////////////////
	
	///////////////////////////////////////////
	//////////////測試嘗試寫入不合法位址//////////////
	///////////////////////////////////////////////
	
	///////////////////1_byte//////////////////////
	#1000 RX = 0;	      //開始02
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////2_byte//////////////////////
	#1000 RX = 0;       //開始 C0(寫入ram[64])1100 0000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////3_byte//////////////////////
	#1000 RX = 0;       //開始 0000_0000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////4_byte//////////////////////
	#1000 RX = 0;       //開始 0000_0000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////5_byte//////////////////////
	#1000 RX = 0;       //開始 0000_0000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////6_byte//////////////////////
	#1000 RX = 0;       //開始 0000_0000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////7_byte//////////////////////
	#1000 RX = 0;       //開始 1100_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////8_byte//////////////////////
	#1000 RX = 0;       //開始 0000_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	#3000 RX = 1;
	
	////////////////////////////////////////////////
	
	///////////////////////////////////////////////
	//////////////再次測試讀出RAM[116]////////////////
	///////////////////////////////////////////////
	
	///////////////////1_byte//////////////////////
	#1000 RX = 0;	      //開始02
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////2_byte//////////////////////
	#1000 RX = 0;       //開始 40(讀出ram[64])0100 0000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////3_byte//////////////////////
	#1000 RX = 0;       //開始 0101_0101
	#1000 RX = 1;       
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////4_byte//////////////////////
	#1000 RX = 0;       //開始 0110_0110
	#1000 RX = 0;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////5_byte//////////////////////
	#1000 RX = 0;       //開始 0111_0111
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	///////////////////6_byte//////////////////////
	#1000 RX = 0;       //開始 1000_1000
	#1000 RX = 0;       
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////7_byte//////////////////////
	#1000 RX = 0;       //開始 1100_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;
	#1000 RX = 1;
	#1000 RX = 1;       //結束
	///////////////////8_byte//////////////////////
	#1000 RX = 0;       //開始 0000_0011
	#1000 RX = 1;       
	#1000 RX = 1;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 0;
	#1000 RX = 1;       //結束
	#3000 RX = 1;
	*/
	////////////////////////////////////////////////
	
	#250000 $stop;      //執行到指定時間後停止
	end
  
	always #10 clk = ~clk;
  
endmodule



